*** SPICE deck for cell Nand{sch} from library Nand
*** Created on Sat Sep 02, 2023 15:24:18
*** Last revised on Sat Sep 02, 2023 17:37:07
*** Written on Sat Sep 02, 2023 17:40:23 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Nand{sch}
Mnmos@0 Out A net@66 gnd NMOS L=0.4U W=2U
Mnmos@1 net@66 B gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd A Out vdd PMOS L=0.4U W=2U
Mpmos@1 vdd B Out vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'Nand{sch}'
vdd vdd 0 DC 1,3
va A 0 pw1 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 pw1 10n 0 20n 5 100n 5 110n 0 
cload out 0 25fF
measure tran tf trig v(out) val=4.5 fall=1 td=4ns trag v(out) val=0.5 fall=1
measure tran tr trig v(out) val=0.5 rais=1 td=4ns trag v(out) val=4.5 rais=1
tran 50n
include C:\Users\soFTech\Downloads\22nm-2.txt
.END
