*** SPICE deck for cell Inv{sch} from library Invertor
*** Created on Sat Aug 26, 2023 23:25:11
*** Last revised on Sun Aug 27, 2023 00:05:27
*** Written on Sun Aug 27, 2023 00:17:52 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

.global gnd vdd

*** TOP LEVEL CELL: Inv{sch}
Mnmos@0 net@7 net@4 gnd gnd SPICE-Model L=0.4U W=2U
Mpmos@0 vdd net@4 net@7 vdd SPICE-Model L=0.4U W=2U

* Spice Code nodes in cell cell 'Inv{sch}'
vdd vdd 0 DC 5
vin in 0 pwl 10n 0 20n 5 50m 5 60n O
cload out 0 250fF
measure tran tf trig v(out) val=4.5 fall=1 td=8ns trag v(out) val=0.5 fall=1
measure tran tr trig v(out) val=0.5 rais=1 td=50ns trag v(out) val=4.5 rais=1
tran 0 0.1 us
include C:\Electric\C5_models.txt
.END
